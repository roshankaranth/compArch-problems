module test;
    integer i;
    wire p;
    reg q;
    parameter n;


    initial begin
        i = 1;
        q = 1;
        p=4;
    end

endmodule